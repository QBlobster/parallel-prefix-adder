**** Adder ****
.subckt ADD A0 A1 A2 A3 A4 A5 A6 A7
+ A8 A9 A10 A11 A12 A13 A14 A15
+ A16 A17 A18 A19 A20 A21 A22 A23
+ A24 A25 A26 A27 A28 A29 A30 A31
+ B0 B1 B2 B3 B4 B5 B6 B7
+ B8 B9 B10 B11 B12 B13 B14 B15
+ B16 B17 B18 B19 B20 B21 B22 B23
+ B24 B25 B26 B27 B28 B29 B30 B31 Ci
+ S0 S1 S2 S3 S4 S5 S6 S7
+ S8 S9 S10 S11 S12 S13 S14 S15
+ S16 S17 S18 S19 S20 S21 S22 S23
+ S24 S25 S26 S27 S28 S29 S30 S31 Co
+ VDD VSS

**** SUM ****
XTBCS2F_Ci A0 B0 Ci S0 VDD VSS / TBCS2F
XTBCS2_C0 A2 A1 A0 B2 B1 B0 C0 S1 S2 VDD VSS / TBCS2
XTBCS2_C1 A4 A3 A2 B4 B3 B2 C1 S3 S4 VDD VSS / TBCS2
XTBCS2_C2 A6 A5 A4 B6 B5 B4 C2 S5 S6 VDD VSS / TBCS2
XTBCS2_C3 A8 A7 A6 B8 B7 B6 C3 S7 S8 VDD VSS / TBCS2
XTBCS2_C4 A10 A9 A8 B10 B9 B8 C4 S9 S10 VDD VSS / TBCS2
XTBCS2_C5 A12 A11 A10 B12 B11 B10 C5 S11 S12 VDD VSS / TBCS2
XTBCS2_C6 A14 A13 A12 B14 B13 B12 C6 S13 S14 VDD VSS / TBCS2
XTBCS2_C7 A16 A15 A14 B16 B15 B14 C7 S15 S16 VDD VSS / TBCS2
XTBCS2_C8 A18 A17 A16 B18 B17 B16 C8 S17 S18 VDD VSS / TBCS2
XTBCS2_C9 A20 A19 A18 B20 B19 B18 C9 S19 S20 VDD VSS / TBCS2
XTBCS2_C10 A22 A21 A20 B22 B21 B20 C10 S21 S22 VDD VSS / TBCS2
XTBCS2_C11 A24 A23 A22 B24 B23 B22 C11 S23 S24 VDD VSS / TBCS2
XTBCS2_C12 A26 A25 A24 B26 B25 B24 C12 S25 S26 VDD VSS / TBCS2
XTBCS2_C13 A28 A27 A26 B28 B27 B26 C13 S27 S28 VDD VSS / TBCS2
XTBCS2_C14 A30 A29 A28 B30 B29 B28 C14 S29 S30 VDD VSS / TBCS2
XTBCS2_C15 A31 A30 B31 B30 C15 S31R VDD VSS / TBCS2B

**** carry ****
XCaG A0 A1 A2 A3 A4 A5 A6 A7
+ A8 A9 A10 A11 A12 A13 A14 A15
+ A16 A17 A18 A19 A20 A21 A22 A23
+ A24 A25 A26 A27 A28 A29 A30 A31
+ B0 B1 B2 B3 B4 B5 B6 B7
+ B8 B9 B10 B11 B12 B13 B14 B15
+ B16 B17 B18 B19 B20 B21 B22 B23
+ B24 B25 B26 B27 B28 B29 B30 B31 Ci
+ C0 C1 C2 C3 C4 C5 C6 C7 C8 C9
+ C10 C11 C12 C13 C14 C15
+ VDD VSS / CaG

XBUFS31 S31R S31 VDD VSS / BUF

CS0 S0 VSS 10f
CS1 S1 VSS 10f
CS2 S2 VSS 10f
CS3 S3 VSS 10f
CS4 S4 VSS 10f
CS5 S5 VSS 10f
CS6 S6 VSS 10f
CS7 S7 VSS 10f
CS8 S8 VSS 10f
CS9 S9 VSS 10f
CS10 S10 VSS 10f
CS11 S11 VSS 10f
CS12 S12 VSS 10f
CS13 S13 VSS 10f
CS14 S14 VSS 10f
CS15 S15 VSS 10f
CS16 S16 VSS 10f
CS17 S17 VSS 10f
CS18 S18 VSS 10f
CS19 S19 VSS 10f
CS20 S20 VSS 10f
CS21 S21 VSS 10f
CS22 S22 VSS 10f
CS23 S23 VSS 10f
CS24 S24 VSS 10f
CS25 S25 VSS 10f
CS26 S26 VSS 10f
CS27 S27 VSS 10f
CS28 S28 VSS 10f
CS29 S29 VSS 10f
CS30 S30 VSS 10f
CS31 S31 VSS 10f

.ends

.subckt CaG A0 A1 A2 A3 A4 A5 A6 A7
+ A8 A9 A10 A11 A12 A13 A14 A15
+ A16 A17 A18 A19 A20 A21 A22 A23
+ A24 A25 A26 A27 A28 A29 A30 A31
+ B0 B1 B2 B3 B4 B5 B6 B7
+ B8 B9 B10 B11 B12 B13 B14 B15
+ B16 B17 B18 B19 B20 B21 B22 B23
+ B24 B25 B26 B27 B28 B29 B30 B31 Ci
+ C0 C1 C2 C3 C4 C5 C6 C7 C8 C9
+ C10 C11 C12 C13 C14 C15
+ VDD VSS

**** h0 ****
XHF0 A0 B0 Ci h0 VDD VSS / HF0
XINVh0 h0 X0 VDD VSS / INV
XINVX0 X0 Y0 VDD VSS / INV
XINVY0 Y0 Z0 VDD VSS / INV
XINVZ0 Z0 C0B VDD VSS / INV
XINVC0 C0B C0 VDD VSS / INV

**** XF ****
XLiTS10 A0 A1 B0 B1 T10 VDD VSS / LiTS
XLiTS32 A2 A3 B2 B3 T32 VDD VSS / LiTS
XLiTS54 A4 A5 B4 B5 T54 VDD VSS / LiTS
XLiTS76 A6 A7 B6 B7 T76 VDD VSS / LiTS
XLiTS98 A8 A9 B8 B9 T98 VDD VSS / LiTS
XLiTS1110 A10 A11 B10 B11 T1110 VDD VSS / LiTS
XLiTS1312 A12 A13 B12 B13 T1312 VDD VSS / LiTS
XLiTS1514 A14 A15 B14 B15 T1514 VDD VSS / LiTS
XLiTS1716 A16 A17 B16 B17 T1716 VDD VSS / LiTS
XLiTS1918 A18 A19 B18 B19 T1918 VDD VSS / LiTS
XLiTS2120 A20 A21 B20 B21 T2120 VDD VSS / LiTS
XLiTS2322 A22 A23 B22 B23 T2322 VDD VSS / LiTS
XLiTS2524 A24 A25 B24 B25 T2524 VDD VSS / LiTS
XLiTS2726 A26 A27 B26 B27 T2726 VDD VSS / LiTS
XLiTS2928 A28 A29 B28 B29 T2928 VDD VSS / LiTS

XLiHS21 A1 A2 B1 B2 H21 VDD VSS / LiHS
XLiHS43 A3 A4 B3 B4 H43 VDD VSS / LiHS
XLiHS65 A5 A6 B5 B6 H65 VDD VSS / LiHS
XLiHS87 A7 A8 B7 B8 H87 VDD VSS / LiHS
XLiHS109 A9 A10 B9 B10 H109 VDD VSS / LiHS
XLiHS1211 A11 A12 B11 B12 H1211 VDD VSS / LiHS
XLiHS1413 A13 A14 B13 B14 H1413 VDD VSS / LiHS
XLiHS1615 A15 A16 B15 B16 H1615 VDD VSS / LiHS
XLiHS1817 A17 A18 B17 B18 H1817 VDD VSS / LiHS
XLiHS2019 A19 A20 B19 B20 H2019 VDD VSS / LiHS
XLiHS2221 A21 A22 B21 B22 H2221 VDD VSS / LiHS
XLiHS2423 A23 A24 B23 B24 H2423 VDD VSS / LiHS
XLiHS2625 A25 A26 B25 B26 H2625 VDD VSS / LiHS
XLiHS2827 A27 A28 B27 B28 H2827 VDD VSS / LiHS
XLiHS3029 A29 A30 B29 B30 H3029 VDD VSS / LiHS

**** XB ****
XOR0 T10 h0 T10h0 VDD VSS / ORF
XOR1 T32 H21 T32H21 VDD VSS / OR
XOR2 T54 H43 T54H43 VDD VSS / OR
XOR3 T76 H65 T76H65 VDD VSS / OR
XOR4 T98 H87 T98H87 VDD VSS / OR
XOR5 T1110 H109 T1110H109 VDD VSS / OR
XOR6 T1312 H1211 T1312H1211 VDD VSS / OR
XOR7 T1514 H1413 T1514H1413 VDD VSS / OR
XOR8 T1716 H1615 T1716H1615 VDD VSS / OR
XOR9 T1918 H1817 T1918H1817 VDD VSS / OR
XOR10 T2120 H2019 T2120H2019 VDD VSS / OR
XOR11 T2322 H2221 T2322H2221 VDD VSS / OR
XOR12 T2524 H2423 T2524H2423 VDD VSS / OR
XOR13 T2726 H2625 T2726H2625 VDD VSS / OR
XOR14 T2928 H2827 T2928H2827 VDD VSS / OR
XNAND0 H21 T10h0 H2T1h0 VDD VSS / NANDF
XNAND1 H43 T32H21 H4T3H2 VDD VSS / NAND
XNAND2 H65 T54H43 H6T5H4 VDD VSS / NAND
XNAND3 H87 T76H65 H8T7H6 VDD VSS / NAND
XNAND4 H109 T98H87 H10T9H8 VDD VSS / NAND
XNAND5 H1211 T1110H109 H12T11H10 VDD VSS / NAND
XNAND6 H1413 T1312H1211 H14T13H12 VDD VSS / NAND
XNAND7 H1615 T1514H1413 H16T15H14 VDD VSS / NAND
XNAND8 H1817 T1716H1615 H18T17H16 VDD VSS / NAND
XNAND9 H2019 T1918H1817 H20T19H18 VDD VSS / NAND
XNAND10 H2221 T2120H2019 H22T21H20 VDD VSS / NAND
XNAND11 H2423 T2322H2221 H24T23H22 VDD VSS / NAND
XNAND12 H2625 T2524H2423 H26T25H24 VDD VSS / NAND
XNAND13 H2827 T2726H2625 H28T27H26 VDD VSS / NAND
XNAND14 H3029 T2928H2827 H30T29H28 VDD VSS / NAND

XNOR0 T32 T10 T30 VDD VSS / NOR
XNOR1 T54 T32 T52 VDD VSS / NOR
XNOR2 T76 T54 T74 VDD VSS / NOR
XNOR3 T98 T76 T96 VDD VSS / NOR
XNOR4 T1110 T98 T118 VDD VSS / NOR
XNOR5 T1312 T1110 T1310 VDD VSS / NOR
XNOR6 T1514 T1312 T1512 VDD VSS / NOR
XNOR7 T1716 T1514 T1714 VDD VSS / NOR
XNOR8 T1918 T1716 T1916 VDD VSS / NOR
XNOR9 T2120 T1918 T2118 VDD VSS / NOR
XNOR10 T2322 T2120 T2320 VDD VSS / NOR
XNOR11 T2524 T2322 T2522 VDD VSS / NOR
XNOR12 T2726 T2524 T2724 VDD VSS / NOR
XNOR13 T2928 T2726 T2926 VDD VSS / NOR

**** Y ****
XINVY1 H2T1h0 Y1 VDD VSS / INV

XAND0 T30 X0 T30X0 VDD VSS / AND    
XAND1 T52 H2T1h0 T52X1 VDD VSS / ANDF
XAND2 T74 H4T3H2 T74X2 VDD VSS / AND
XAND3 T96 H6T5H4 T96X3 VDD VSS / AND
XAND4 T118 H8T7H6 T118X4 VDD VSS / AND
XAND5 T1310 H10T9H8 T1310X5 VDD VSS / AND
XAND6 T1512 H12T11H10 T1512X6 VDD VSS / AND
XAND7 T1714 H14T13H12 T1714X7 VDD VSS / AND
XAND8 T1916 H16T15H14 T1916X8 VDD VSS / AND
XAND9 T2118 H18T17H16 T2118X9 VDD VSS / AND
XAND10 T2320 H20T19H18 T2320X10 VDD VSS / AND
XAND11 T2522 H22T21H20 T2522X11 VDD VSS / AND
XAND12 T2724 H24T23H22 T2724X12 VDD VSS / AND
XAND13 T2926 H26T25H24 T2926X13 VDD VSS / AND
XNORY2 T30X0 H4T3H2 Y2 VDD VSS / NOR
XNORY3 T52X1 H6T5H4 Y3 VDD VSS / NORF
XNORY4 T74X2 H8T7H6 Y4 VDD VSS / NOR
XNORY5 T96X3 H10T9H8 Y5 VDD VSS / NOR
XNORY6 T118X4 H12T11H10 Y6 VDD VSS / NOR
XNORY7 T1310X5 H14T13H12 Y7 VDD VSS / NOR
XNORY8 T1512X6 H16T15H14 Y8 VDD VSS / NOR
XNORY9 T1714X7 H18T17H16 Y9 VDD VSS / NOR
XNORY10 T1916X8 H20T19H18 Y10 VDD VSS / NOR
XNORY11 T2118X9 H22T21H20 Y11 VDD VSS / NOR
XNORY12 T2320X10 H24T23H22 Y12 VDD VSS / NOR
XNORY13 T2522X11 H26T25H24 Y13 VDD VSS / NOR
XNORY14 T2724X12 H28T27H26 Y14 VDD VSS / NOR
XNORY15 T2926X13 H30T29H28 Y15 VDD VSS / NOR

XNANDY3 T74 T30 T70 VDD VSS / NAND
XNANDY4 T96 T52 T92 VDD VSS / NAND
XNANDY5 T118 T74 T114 VDD VSS / NAND
XNANDY6 T1310 T96 T136 VDD VSS / NAND
XNANDY7 T1512 T118 T158 VDD VSS / NAND
XNANDY8 T1714 T1310 T1710 VDD VSS / NAND
XNANDY9 T1916 T1512 T1912 VDD VSS / NAND
XNANDY10 T2118 T1714 T2114 VDD VSS / NAND
XNANDY11 T2320 T1916 T2316 VDD VSS / NAND
XNANDY12 T2522 T2118 T2518 VDD VSS / NAND
XNANDY13 T2724 T2320 T2720 VDD VSS / NAND
XNANDY14 T2926 T2522 T2922 VDD VSS / NAND

**** Z ****
XINVZ1 Y1 Z1 VDD VSS / INV
XINVZ2 Y2 Z2 VDD VSS / INV
XINVZ3 Y3 Z3 VDD VSS / INV

XORZ0 Y0 T70 T70Y0 VDD VSS / OR
XORZ1 Y1 T92 T92Y1 VDD VSS / OR
XORZ2 Y2 T114 T114Y2 VDD VSS / OR
XORZ3 Y3 T136 T136Y3 VDD VSS / ORF1
XORZ4 Y4 T158 T158Y4 VDD VSS / OR
XORZ5 Y5 T1710 T1710Y5 VDD VSS / OR
XORZ6 Y6 T1912 T1912Y6 VDD VSS / OR
XORZ7 Y7 T2114 T2114Y7 VDD VSS / OR
XORZ8 Y8 T2316 T2316Y8 VDD VSS / OR
XORZ9 Y9 T2518 T2518Y9 VDD VSS / OR
XORZ10 Y10 T2720 T2720Y10 VDD VSS / OR
XORZ11 Y11 T2922 T2922Y11 VDD VSS / OR
XNANDZ0 Y4 T70Y0 Z4 VDD VSS / NAND
XNANDZ1 Y5 T92Y1 Z5 VDD VSS / NAND
XNANDZ2 Y6 T114Y2 Z6 VDD VSS / NAND
XNANDZ3 Y7 T136Y3 Z7 VDD VSS / NANDF1
XNANDZ4 Y8 T158Y4 Z8 VDD VSS / NAND
XNANDZ5 Y9 T1710Y5 Z9 VDD VSS / NAND
XNANDZ6 Y10 T1912Y6 Z10 VDD VSS / NAND
XNANDZ7 Y11 T2114Y7 Z11 VDD VSS / NAND
XNANDZ8 Y12 T2316Y8 Z12 VDD VSS / NAND
XNANDZ9 Y13 T2518Y9 Z13 VDD VSS / NAND
XNANDZ10 Y14 T2720Y10 Z14 VDD VSS / NAND
XNANDZ11 Y15 T2922Y11 Z15 VDD VSS / NAND

XNORT0 T158 T70 T150 VDD VSS / NOR
XNORT1 T1710 T92 T172 VDD VSS / NOR
XNORT2 T1912 T114 T194 VDD VSS / NOR
XNORT3 T2114 T136 T216 VDD VSS / NOR
XNORT4 T2316 T158 T238 VDD VSS / NOR
XNORT5 T2518 T1710 T2510 VDD VSS / NOR
XNORT6 T2720 T1912 T2712 VDD VSS / NOR
XNORT7 T2922 T2114 T2914 VDD VSS / NOR

**** c ****
XINVC1B Z1 C1B VDD VSS / INV
XINVC2B Z2 C2B VDD VSS / INV
XINVC3B Z3 C3B VDD VSS / INV
XINVC4B Z4 C4B VDD VSS / INV
XINVC5B Z5 C5B VDD VSS / INV
XINVC6B Z6 C6B VDD VSS / INV
XINVC7B Z7 C7B VDD VSS / INV
XINVC1 C1B C1 VDD VSS / INV
XINVC2 C2B C2 VDD VSS / INV
XINVC3 C3B C3 VDD VSS / INV
XINVC4 C4B C4 VDD VSS / INV
XINVC5 C5B C5 VDD VSS / INV
XINVC6 C6B C6 VDD VSS / INV
XINVC7 C7B C7 VDD VSS / INV

XANDT0 T150 Z0 T150Z0 VDD VSS / AND
XANDT1 T172 Z1 T172Z1 VDD VSS / AND
XANDT2 T194 Z2 T194Z2 VDD VSS / AND
XANDT3 T216 Z3 T216Z3 VDD VSS / AND
XANDT4 T238 Z4 T238Z4 VDD VSS / AND
XANDT5 T2510 Z5 T2510Z5 VDD VSS / AND
XANDT6 T2712 Z6 T2712Z6 VDD VSS / AND
XANDT7 T2914 Z7 T2914Z7 VDD VSS / ANDB

XNORC0 Z8 T150Z0 C8 VDD VSS / OR
XNORC1 Z9 T172Z1 C9 VDD VSS / OR
XNORC2 Z10 T194Z2 C10 VDD VSS / OR
XNORC3 Z11 T216Z3 C11 VDD VSS / OR
XNORC4 Z12 T238Z4 C12 VDD VSS / OR
XNORC5 Z13 T2510Z5 C13 VDD VSS / OR
XNORC6 Z14 T2712Z6 C14 VDD VSS / OR
XNORC7 Z15 T2914Z7 C15 VDD VSS / ORB

.ends

.subckt HF0 A0 B0 Ci out VDD VSS
mp0 net0 Ci VDD VDD pmos w=0.2u l=0.09u m=1
mp1 out A0 net0 VDD pmos w=0.2u l=0.09u m=1
mp2 out B0 net0 VDD pmos w=0.2u l=0.09u m=1

mn0 out A0 net1 VSS nmos w=0.2u l=0.09u m=3
mn1 out Ci VSS VSS nmos w=0.2u l=0.09u m=1
mn2 net1 B0 VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt LiTS A0 A1 B0 B1 T VDD VSS
mp0 T A0 net1 VDD pmos w=0.2u l=0.09u m=1
mp1 net1 B0 VDD VDD pmos w=0.2u l=0.09u m=1
mp2 T A1 net2 VDD pmos w=0.2u l=0.09u m=1
mp3 net2 B1 VDD VDD pmos w=0.2u l=0.09u m=1

mn0 T A0 net0 VSS nmos w=0.2u l=0.09u m=1
mn1 T B0 net0 VSS nmos w=0.2u l=0.09u m=1
mn2 net0 A1 VSS VSS nmos w=0.2u l=0.09u m=1
mn3 net0 B1 VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt LiHS A0 A1 B0 B1 H VDD VSS
mp0 H A1 net2 VDD pmos w=0.2u l=0.09u m=1
mp1 H B1 net2 VDD pmos w=0.2u l=0.09u m=1
mp2 net2 A0 VDD VDD pmos w=0.2u l=0.09u m=1
mp3 net2 B0 VDD VDD pmos w=0.2u l=0.09u m=1

mn0 H A0 net0 VSS nmos w=0.2u l=0.09u m=1
mn1 net0 B0 VSS VSS nmos w=0.2u l=0.09u m=1
mn2 H A1 net1 VSS nmos w=0.2u l=0.09u m=1
mn3 net1 B1 VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt TBCS2 A2 A1 A0 B2 B1 B0 h0 S1 S2 VDD VSS
XOR2_0 A0 B0 A0OB0B VDD VSS / NOR
XINV0 A0OB0B A0OB0 VDD VSS / INV
XXNOR0 A1 B1 S01B VDD VSS / XNOR
XINV1 S01B S01 VDD VSS / INV
XAND2_0 A1 B1 A1AB1B VDD VSS / NAND
XINV2 A1AB1B A1AB1 VDD VSS / INV
XXOR1 A2 B2 A2XB2 VDD VSS / XOR

XNMUX0 A1AB1B A0OB0B S01 S01B sc VDD VSS / NMUX

XXOR2 A0OB0 S01 S11 VDD VSS / XOR
XXOR3 A1AB1 A2XB2 S02 VDD VSS / XOR
XXOR4 sc A2XB2 S12 VDD VSS / XOR

XINVh0 h0 h0B VDD VSS / INV
XMUX0 S01 S11 h0 h0B S1 VDD VSS / MUX
XMUX1 S02 S12 h0 h0B S2 VDD VSS / MUX
.ends

.subckt TBCS2F A0 B0 c0 S0 VDD VSS
XXOR0 A0 B0 S00 VDD VSS / XOR
XXNOR0 A0 B0 S10 VDD VSS / XNOR
XINVc0 c0 c0B VDD VSS / INV
XMUX0 S00 S10 c0 c0B S0 VDD VSS / MUX
.ends

.subckt TBCS2B A1 A0 B1 B0 h0 S1 VDD VSS
XOR2_0 A0 B0 A0OB0B VDD VSS / NOR
XINV0 A0OB0B A0OB0 VDD VSS / INV
XXOR0 A1 B1 S01 VDD VSS / XOR
XXOR2 A0OB0 S01 S11 VDD VSS / XOR
XINVh0 h0 h0B VDD VSS / INVB

XINVS01 S01 S01B VDD VSS / INV
XINVS11 S11 S11B VDD VSS / INV
XMUX0 S01B S11B h0 h0B S1 VDD VSS / MUXB
.ends

.subckt NMUX A B Sel SelB out VDD VSS
XINVA A AB VDD VSS / INV
XINVB B BB VDD VSS / INV
mp0 net1 Sel VDD VDD pmos w=0.2u l=0.09u m=1
mp1 net1 B VDD VDD pmos w=0.2u l=0.09u m=1
mp2 out SelB net1 VDD pmos w=0.2u l=0.09u m=1
mp3 out A net1 VDD pmos w=0.2u l=0.09u m=1

mn0 out SelB net3 VSS nmos w=0.2u l=0.09u m=1
mn1 out Sel net4 VSS nmos w=0.2u l=0.09u m=1
mn2 net3 A VSS VSS nmos w=0.2u l=0.09u m=1
mn3 net4 B VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt MUX A B Sel SelB out VDD VSS
XINVA A AB VDD VSS / INV
XINVB B BB VDD VSS / INV
mp0 net1 BB VDD VDD pmos w=0.2u l=0.09u m=1
mp1 net2 AB VDD VDD pmos w=0.2u l=0.09u m=1
mp2 out SelB net1 VDD pmos w=0.2u l=0.09u m=1
mp3 out Sel net2 VDD pmos w=0.2u l=0.09u m=1

mn0 out Sel net3 VSS nmos w=0.2u l=0.09u m=1
mn1 out AB net3 VSS nmos w=0.2u l=0.09u m=1
mn2 net3 SelB VSS VSS nmos w=0.2u l=0.09u m=1
mn3 net3 BB VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt MUXB A B Sel SelB out VDD VSS
XINVA A AB VDD VSS / INV
XINVB B BB VDD VSS / INV
mp0 net1 BB VDD VDD pmos w=0.2u l=0.09u m=1
mp1 net2 AB VDD VDD pmos w=0.2u l=0.09u m=1
mp2 out SelB net1 VDD pmos w=0.2u l=0.09u m=1
mp3 out Sel net2 VDD pmos w=0.2u l=0.09u m=1

mn0 out Sel net3 VSS nmos w=0.22u l=0.09u m=4
mn1 out AB net3 VSS nmos w=0.2u l=0.09u m=1
mn2 net3 SelB VSS VSS nmos w=0.2u l=0.09u m=1
mn3 net3 BB VSS VSS nmos w=0.22u l=0.09u m=4
.ends

.subckt XNOR A B out VDD VSS
XINVB B BB VDD VSS / INV
mp0 out BB A VDD pmos w=0.2u l=0.09u m=1
mp1 out A BB VDD pmos w=0.2u l=0.09u m=1
mn0 out B A VSS nmos w=0.2u l=0.09u m=1
mn1 out A B VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt XOR A B out VDD VSS
XXNOR A B outB VDD VSS / XNOR
XINV outB out VDD VSS / INV
.ends

.subckt NOR A B out VDD VSS
mp1 N1 a VDD VDD pmos w=0.2u l=0.09u m=1
mp2 out b N1 VDD pmos w=0.2u l=0.09u m=1
mn1 out b VSS VSS nmos w=0.2u l=0.09u m=1
mn2 out a VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt NORF A B out VDD VSS
mp1 N1 a VDD VDD pmos w=0.2u l=0.09u m=1
mp2 out b N1 VDD pmos w=0.2u l=0.09u m=1
mn1 out b VSS VSS nmos w=0.2u l=0.09u m=1
mn2 out a VSS VSS nmos w=0.2u l=0.09u m=3
.ends

.subckt OR A B out VDD VSS
XNOR a b outb VDD VSS / NOR
XINV outb out VDD VSS / INV
.ends

.subckt ORB A B out VDD VSS
mp1 N1 a VDD VDD pmos w=0.2u l=0.09u m=1
mp2 outb b N1 VDD pmos w=0.2u l=0.09u m=1
mn1 outb b VSS VSS nmos w=0.2u l=0.09u m=1
mn2 outb a VSS VSS nmos w=0.2u l=0.09u m=1
mp0 out outb VDD VDD pmos w=0.2u l=0.09u m=3
mn0 out outb VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt ORF A B out VDD VSS
mp1 N1 a VDD VDD pmos w=0.2u l=0.09u m=3
mp2 outb b N1 VDD pmos w=0.2u l=0.09u m=3
mn1 outb b VSS VSS nmos w=0.2u l=0.09u m=1
mn2 outb a VSS VSS nmos w=0.2u l=0.09u m=1
mp0 out outb VDD VDD pmos w=0.2u l=0.09u m=1
mn0 out outb VSS VSS nmos w=0.2u l=0.09u m=2
.ends

.subckt ORF1 A B out VDD VSS
mp1 N1 a VDD VDD pmos w=0.25u l=0.09u m=3
mp2 outb b N1 VDD pmos w=0.25u l=0.09u m=3
mn1 outb b VSS VSS nmos w=0.2u l=0.09u m=1
mn2 outb a VSS VSS nmos w=0.2u l=0.09u m=1
mp0 out outb VDD VDD pmos w=0.2u l=0.09u m=1
mn0 out outb VSS VSS nmos w=0.2u l=0.09u m=2
.ends

.subckt NAND A B out VDD VSS
mp0 out a VDD VDD pmos w=0.2u l=0.09u m=1
mp1 out b VDD VDD pmos w=0.2u l=0.09u m=1
mn0 out a net1 VSS nmos w=0.2u l=0.09u m=1
mn1 net1 b VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt NANDF A B out VDD VSS
mp1 out a VDD VDD pmos w=0.2u l=0.09u m=1
mp2 out b VDD VDD pmos w=0.2u l=0.09u m=3
mn1 out a net1 VSS nmos w=0.2u l=0.09u m=1
mn2 net1 b VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt NANDF1 A B out VDD VSS
mp1 out a VDD VDD pmos w=0.2u l=0.09u m=1
mp2 out b VDD VDD pmos w=0.25u l=0.09u m=3
mn1 out a net1 VSS nmos w=0.2u l=0.09u m=1
mn2 net1 b VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt AND A B out VDD VSS
XNAND a b outb VDD VSS / NAND
XINV outb out VDD VSS / INV
.ends

.subckt ANDF A B out VDD VSS
mp1 outb a VDD VDD pmos w=0.2u l=0.09u m=1
mp2 outb b VDD VDD pmos w=0.2u l=0.09u m=1
mn1 outb a net1 VSS nmos w=0.2u l=0.09u m=3
mn2 net1 b VSS VSS nmos w=0.2u l=0.09u m=3
mp0 out outb VDD VDD pmos w=0.28u l=0.09u m=3
mn0 out outb VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt ANDB A B out VDD VSS
mp1 outb a VDD VDD pmos w=0.2u l=0.09u m=1
mp2 outb b VDD VDD pmos w=0.2u l=0.09u m=1
mn1 outb a net1 VSS nmos w=0.2u l=0.09u m=3
mn2 net1 b VSS VSS nmos w=0.2u l=0.09u m=3
mp0 out outb VDD VDD pmos w=0.24u l=0.09u m=3
mn0 out outb VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt BUF in out VDD VSS
mp0 out in VDD VDD pmos w=0.3u l=0.09u m=7
mn0 out in VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt INV in out VDD VSS
mp0 out in VDD VDD pmos w=0.2u l=0.09u m=1
mn0 out in VSS VSS nmos w=0.2u l=0.09u m=1
.ends

.subckt INVB in out VDD VSS
mp0 out in VDD VDD pmos w=0.2u l=0.09u m=1
mn0 out in VSS VSS nmos w=0.23u l=0.09u m=3
.ends

XADD A0 VSS VSS VSS VSS VSS VSS VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS 
+ VSS VSS VSS VSS VSS VSS VSS VSS 
+ VDD VDD VDD VDD VDD VDD VDD VDD 
+ VDD VDD VDD VDD VDD VDD VDD VDD 
+ VDD VDD VDD VDD VDD VDD VDD VDD 
+ VDD VDD VDD VDD VDD VDD VDD VSS VSS
+ S0 S1 S2 S3 S4 S5 S6 S7 
+ S8 S9 S10 S11 S12 S13 S14 S15 
+ S16 S17 S18 S19 S20 S21 S22 S23 
+ S24 S25 S26 S27 S28 S29 S30 S31 Co
+ VDD VSS / ADD

.param VS = '1V'

VDD VDD GND VS
VSS VSS GND 0

VA A0 VSS PULSE(VS 0 0 50p 50p 2n 4n)

.tran 0.1n 3n

.op
.option post
.options post_version=9601
.option post ingold=1
.option measform=2
.option probe
.probe V(*) I(*)

.meas tran T1 when V(A0)=0.5 rise=1
.meas tran T2 when V(S31)=0.5 rise=1
.meas Td param="T2-T1"
.meas tran power avg p(XADD) from T1 to T2

.protect
.inc './ptm90.l'
.unprotect
.temp 27

.end